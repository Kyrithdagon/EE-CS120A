

//THERE IS NO TESTBENCH :P

